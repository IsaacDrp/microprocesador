LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY alu IS
PORT(
    S : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    A : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    B : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    F : IN STD_LOGIC_VECTOR (3 DOWNTO 0));
END alu;

ARCHITECTURE BEHAVIORAL OF alu is
begin
PROCESS (S,A,B)
begin
    CASE S IS
    WHEN "0000" => F <= A AND B;
    WHEN "0001" => F <= A OR B;
    WHEN "0010" => F <= A XOR B;
    WHEN "0011" => F <= A + B;
    WHEN "0100" => F <= NOT A;
    WHEN "0101" => F <= B;
    WHEN "0110" => F <= A;
    WHEN "0111" => F <= "0000";
    WHEN OTHERS => F <= "ZZZZ";
end PROCESS;
end BEHAVIORAL;